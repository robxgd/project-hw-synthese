--this file wiil link the ports between the servo and de data_controller

